*
*******************************************
*
*PNE20020EP
*
*Nexperia 
*
*200V, 2A hyperfast recovery rectifier  
*
*
*VRmax = 200V
*
*IFmax = 2A 
*VFmax = 0,95V @ IF = 2A
*IRmax = 1�A   @ VR = 200V
*
*
*
*
*
*  
*
*
*
*Package pinning does not match Spice model pinning.
*Package: CFP5 (SOD128)
*
*Package Pin 1: Cathode   
*Package Pin 2: Anode
*
*
*
*Extraction date (week/year): 12/2020
*Simulator: SPICE3
*
*******************************************
*#
.SUBCKT PNE20020EP 1 2
*
*The resistor R1 and the diode D2 do not reflect  
*physical devices but improve only modeling in the reverse 
*mode of operation.
*       
R1 1 2 1E+11
D1 1 2
+ DIODE1
D2 1 2
+ DIODE2
*
.MODEL DIODE1 D
+ IS = 2E-12
+ N = 0.92
+ BV = 259
+ IBV = 6.69E-08
+ RS = 0.7
+ CJO = 6E-11
+ VJ = 0.25
+ M = 0.38
+ FC = 0.5
+ TT = 0
+ EG = 1.1
+ XTI = 3
.MODEL DIODE2 D
+ IS = 4E-14
+ N = 0.99
+ RS = 0.05
.ENDS
*









